* Universal Opamp SPICE Macromodels
* Version: v1.1
* Date: 2019-11-23
* 
* Written in 2019 by Ste Kulov, HD Retrovision LLC.
* Later modified by KiCad developers
* To the extent possible under law, the author(s) have dedicated all copyright
* and related and neighboring rights to this software to the public domain worldwide. 
* This software is distributed without any warranty. 
* You should have received a copy of the CC0 Public Domain Dedication along with this software.
* If not, see <http://creativecommons.org/publicdomain/zero/1.0/>.
* 
*****************************************
*************
* CHANGELOG *
*************
* ---------------------------------------
* v1.0
* 2019-11-08
* ---------------------------------------
* 1.) Initial Release
* ---------------------------------------
* 
* 
* ---------------------------------------
* v1.1
* 2019-11-23
* ---------------------------------------
* 1.) lvl2:	Removed SW model and replaced all instances with semiconductor diodes.
* 2.) lvl2: Added offsets to the voltage sources to compensate for the new semiconductor junctions.
* ---------------------------------------
* v1.2
* 2022-08-23
* ---------------------------------------
* 1.) Added dual and quad channel models for both lvl1 and lvl2
*****************************************


*****************************************
.subckt uopamp_lvl1 +IN -IN OUT
* Universal Opamp Level 1
* Single pole opamp without voltage rails and referenced to GND
* 
* PINOUT ORDER  1   2   3
* PINOUT ORDER +IN -IN OUT
* 
* Parameters:
* Avol => open-loop voltage gain (V/V), default=100k
* GBW => gain-bandwidth product (Hz), default=100meg
* Rin => differential input resistance (ohm), default=100g
* Rout => open-loop output resistance (ohm), default=1
* 
R1 +IN -IN {Rin}
G1 0 OUT +IN -IN {Avol/Rout}
R2 OUT 0 100g
C3 OUT 0 {Avol/(2*pi*GBW*Rout)}
.param Avol=100k
.param GBW=100meg
.param Rin=100g
.param Rout=1
.param pi=3.1415926535898
.ends

*****************************************
.subckt uopamp_lvl1_2x +IN1 -IN1 OUT1 +IN2 -IN2 OUT2
X1 +IN1 -IN1 OUT1 uopamp_lvl1
X2 +IN2 -IN2 OUT2 uopamp_lvl1
.ends
*****************************************

*****************************************
.subckt uopamp_lvl1_4x +IN1 -IN1 OUT1 +IN2 -IN2 OUT2 +IN3 -IN3 OUT3 +IN4 -IN4 OUT4
X1 +IN1 -IN1 OUT1 uopamp_lvl1 
X2 +IN2 -IN2 OUT2 uopamp_lvl1 
X3 +IN3 -IN3 OUT3 uopamp_lvl1 
X4 +IN4 -IN4 OUT4 uopamp_lvl1 
.ends
*****************************************


*****************************************
.subckt uopamp_lvl2 +IN -IN VCC VEE OUT
* Universal Opamp Level 2
* Single pole opamp with rail saturation, current consumption, current limiting, and input offset voltage
* 
* PINOUT ORDER  1   2   3   4   5
* PINOUT ORDER +IN -IN VCC VEE OUT
* 
* Parameters:
* Avol => open-loop voltage gain (V/V), default=100k
* GBW => gain-bandwidth product (Hz), default=100meg
* Rin => differential input resistance (ohm), default=100g
* Rout => open-loop output resistance (ohm), default=1
* Iq => quiescent supply current (A), default=1m
* Ilimit => maximum output current (A), default=1
* Vrail => voltage between output saturation and each rail (V), default=0
* Vos => input offset voltage (V), default=0
* Vmax => total maximum supply voltage between rails (V), default=50
* 
G1 VCC N001 N002 -IN 1u
G2 VEE N001 N002 -IN 1u
R1 VCC N001 {Avol/1u}
R2 N001 VEE {Avol/1u}
G3 OUT VCC VCC N001 {1/(2*Rout)}
G4 VEE OUT N001 VEE {1/(2*Rout)}
R4 VCC OUT {2*Rout}
R5 OUT VEE {2*Rout}
C1 VCC N001 {1u/(2*pi*GBW)}
C2 N001 VEE {1u/(2*pi*GBW)}
G6 N005 VEE N001 OUT {1/(2*Rout)}
G5 N006 VEE OUT N001 {1/(2*Rout)}
R8 -IN +IN {Rin}
V6 VCC N003 {Vrail+545m}
V7 N008 VEE {Vrail+545m}
V8 N002 +IN {Vos}
V9 OUT N007 {Ilimit-545m}
V10 N004 OUT {Ilimit-545m}
D1 N001 N003 diode
D2 N008 N001 diode
D3 VCC N005 diode
D4 VCC N006 diode
D5 VEE N005 zener
D6 VEE N006 zener
D7 N001 N004 diode
D8 N007 N001 diode
I1 VCC VEE {Iq}
.param Avol = 100k
.param GBW = 100meg
.param Rin = 100g
.param Rout = 1
.param Iq = 1m
.param Ilimit = 1
.param Vrail = 0
.param Vos = 0
.param Vmax = 50
.model diode D(Is=1e-14)
.model zener D(Is=1e-14 BV={Vmax})
.param pi=3.1415926535898
.ends
*****************************************

*****************************************
.subckt uopamp_lvl2_2x VCC VEE +IN1 -IN1 OUT1 +IN2 -IN2 OUT2
X1 +IN1 -IN1 VCC VEE OUT1 uopamp_lvl2 
X2 +IN2 -IN2 VCC VEE OUT2 uopamp_lvl2 
.ends
*****************************************

*****************************************
.subckt uopamp_lvl2_4x VCC VEE +IN1 -IN1 OUT1 +IN2 -IN2 OUT2 +IN3 -IN3 OUT3 +IN4 -IN4 OUT4
X1 +IN1 -IN1 VCC VEE OUT1 uopamp_lvl2 
X2 +IN2 -IN2 VCC VEE OUT2 uopamp_lvl2 
X3 +IN3 -IN3 VCC VEE OUT3 uopamp_lvl2 
X4 +IN4 -IN4 VCC VEE OUT4 uopamp_lvl2 
.ends
*****************************************
